module pl_instmem (a,inst);
    input  [31:0] a;
    output [31:0] inst;
    wire   [31:0] rom [0:31];                                 // (pc)
    assign rom[5'h00] = 32'b00000001000000000000000010010011; // (00)addi x1, x0, 16   x1=00000010
    assign rom[5'h01] = 32'b00000100000000001000001000010011; // (04)addi  x4, x1, 64  x4=00000050
    assign rom[5'h02] = 32'b00000000000000100010010010000011; // (08)lw  x9, 0 (x4)    x9=memory[x4]=000000f2 
    assign rom[5'h03] = 32'b01000000010001001000010000110011; // (0c)sub x8 , x9, x4   x8=x9-x4=000000a2 
    assign rom[5'h04] = 32'b00000000000000001000011001100011; // (10)beq x1, x0, address+12
    assign rom[5'h05] = 32'b00000000000000000000000000000000; // (14)nop
    assign rom[5'h06] = 32'b00000000101000000000000100010011; // (18)addi x2, x0, 10   x2=0000000a
    assign rom[5'h07] = 32'b00000001010000000000000110010011; // (1c)addi x3, x0, 20   x3=00000014
    assign rom[5'h08] = 32'b00000000000000001001011001100011; // (20)bne x1, x0, address+12
    assign rom[5'h09] = 32'b00000000000000000000000000000000; // (24)nop
    assign rom[5'h0a] = 32'b00000000101000000000001010010011; // (28)addi x5, x0, 10   x5=0000000a
    assign rom[5'h0b] = 32'b00000001010000000000001100010011; // (2c)addi x6, x0, 20   x6=00000014
    assign inst = rom[a[6:2]];
endmodule
